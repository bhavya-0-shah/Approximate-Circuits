module BIT_G(output BG, input A, B);

   and (BG, A, B);

endmodule