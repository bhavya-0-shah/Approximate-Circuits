module BIT_P(output BP, input A, B);

   xor (BP, A, B);

endmodule